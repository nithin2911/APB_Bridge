package my_package;
 	`include "uvm_macros.svh"
   	import uvm_pkg::*;
	`include "my_test.svh"
endpackage
